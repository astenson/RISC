`include "multBlock.v"

module mult();
  wire zero = 1'b0;
  wire [15:0] carry0, carry1, carry2, carry3, carry4, carry5, carry6, carry7, carry8, carry9, carry10, carry11, carry12, carry13, carry14, carry15;
  wire [14:0] add0, add1, add2, add3, add4, add5, add6, add7, add8, add9, add10, add11, add12, add13, add14, add15;
  reg [15:0] A = 16'b0000_0000_0000_0010;
  reg [15:0] B = 16'b0000_0000_0000_0010;
  wire [31:0] result;
  //1st row of multiplier blocks
  multBlock mult00(.x(A[0]),.y(zero),.alt(B[0]),.Cin(zero),.S(result[0]),.Cout(carry0[0]));
  multBlock mult01(.x(A[1]),.y(zero),.alt(B[0]),.Cin(carry0[0]),.S(add0[0]),.Cout(carry0[1]));
  multBlock mult02(.x(A[2]),.y(zero),.alt(B[0]),.Cin(carry0[1]),.S(add0[1]),.Cout(carry0[2]));
  multBlock mult03(.x(A[3]),.y(zero),.alt(B[0]),.Cin(carry0[2]),.S(add0[2]),.Cout(carry0[3]));
  multBlock mult04(.x(A[4]),.y(zero),.alt(B[0]),.Cin(carry0[3]),.S(add0[3]),.Cout(carry0[4]));
  multBlock mult05(.x(A[5]),.y(zero),.alt(B[0]),.Cin(carry0[4]),.S(add0[4]),.Cout(carry0[5]));
  multBlock mult06(.x(A[6]),.y(zero),.alt(B[0]),.Cin(carry0[5]),.S(add0[5]),.Cout(carry0[6]));
  multBlock mult07(.x(A[7]),.y(zero),.alt(B[0]),.Cin(carry0[6]),.S(add0[6]),.Cout(carry0[7]));
  multBlock mult08(.x(A[8]),.y(zero),.alt(B[0]),.Cin(carry0[7]),.S(add0[7]),.Cout(carry0[8]));
  multBlock mult09(.x(A[9]),.y(zero),.alt(B[0]),.Cin(carry0[8]),.S(add0[8]),.Cout(carry0[9]));
  multBlock mult010(.x(A[10]),.y(zero),.alt(B[0]),.Cin(carry0[9]),.S(add0[9]),.Cout(carry0[10]));
  multBlock mult011(.x(A[11]),.y(zero),.alt(B[0]),.Cin(carry0[10]),.S(add0[10]),.Cout(carry0[11]));
  multBlock mult012(.x(A[12]),.y(zero),.alt(B[0]),.Cin(carry0[11]),.S(add0[11]),.Cout(carry0[12]));
  multBlock mult013(.x(A[13]),.y(zero),.alt(B[0]),.Cin(carry0[12]),.S(add0[12]),.Cout(carry0[13]));
  multBlock mult014(.x(A[14]),.y(zero),.alt(B[0]),.Cin(carry0[13]),.S(add0[13]),.Cout(carry0[14]));
  multBlock mult015(.x(A[15]),.y(zero),.alt(B[0]),.Cin(carry0[14]),.S(add0[14]),.Cout(carry0[15]));
  //2nd row of multiplier blocks
  multBlock mult10(.x(A[0]),.y(add0[0]),.alt(B[1]),.Cin(zero),.S(result[1]),.Cout(carry1[0]));
  multBlock mult11(.x(A[1]),.y(add0[1]),.alt(B[1]),.Cin(carry1[0]),.S(add1[0]),.Cout(carry1[1]));
  multBlock mult12(.x(A[2]),.y(add0[2]),.alt(B[1]),.Cin(carry1[1]),.S(add1[1]),.Cout(carry1[2]));
  multBlock mult13(.x(A[3]),.y(add0[3]),.alt(B[1]),.Cin(carry1[2]),.S(add1[2]),.Cout(carry1[3]));
  multBlock mult14(.x(A[4]),.y(add0[4]),.alt(B[1]),.Cin(carry1[3]),.S(add1[3]),.Cout(carry1[4]));
  multBlock mult15(.x(A[5]),.y(add0[5]),.alt(B[1]),.Cin(carry1[4]),.S(add1[4]),.Cout(carry1[5]));
  multBlock mult16(.x(A[6]),.y(add0[6]),.alt(B[1]),.Cin(carry1[5]),.S(add1[5]),.Cout(carry1[6]));
  multBlock mult17(.x(A[7]),.y(add0[7]),.alt(B[1]),.Cin(carry1[6]),.S(add1[6]),.Cout(carry1[7]));
  multBlock mult18(.x(A[8]),.y(add0[8]),.alt(B[1]),.Cin(carry1[7]),.S(add1[7]),.Cout(carry1[8]));
  multBlock mult19(.x(A[9]),.y(add0[9]),.alt(B[1]),.Cin(carry1[8]),.S(add1[8]),.Cout(carry1[9]));
  multBlock mult110(.x(A[10]),.y(add0[10]),.alt(B[1]),.Cin(carry1[9]),.S(add1[9]),.Cout(carry1[10]));
  multBlock mult111(.x(A[11]),.y(add0[11]),.alt(B[1]),.Cin(carry1[10]),.S(add1[10]),.Cout(carry1[11]));
  multBlock mult112(.x(A[12]),.y(add0[12]),.alt(B[1]),.Cin(carry1[11]),.S(add1[11]),.Cout(carry1[12]));
  multBlock mult113(.x(A[13]),.y(add0[13]),.alt(B[1]),.Cin(carry1[12]),.S(add1[12]),.Cout(carry1[13]));
  multBlock mult114(.x(A[14]),.y(add0[14]),.alt(B[1]),.Cin(carry1[13]),.S(add1[13]),.Cout(carry1[14]));
  multBlock mult115(.x(A[15]),.y(carry0[15]),.alt(B[1]),.Cin(carry1[14]),.S(add1[14]),.Cout(carry1[15]));
  //3rd row of multiplier blocks
  multBlock mult20(.x(A[0]),.y(add1[0]),.alt(B[2]),.Cin(zero),.S(result[2]),.Cout(carry2[0]));
  multBlock mult21(.x(A[1]),.y(add1[1]),.alt(B[2]),.Cin(carry2[0]),.S(add2[0]),.Cout(carry2[1]));
  multBlock mult22(.x(A[2]),.y(add1[2]),.alt(B[2]),.Cin(carry2[1]),.S(add2[1]),.Cout(carry2[2]));
  multBlock mult23(.x(A[3]),.y(add1[3]),.alt(B[2]),.Cin(carry2[2]),.S(add2[2]),.Cout(carry2[3]));
  multBlock mult24(.x(A[4]),.y(add1[4]),.alt(B[2]),.Cin(carry2[3]),.S(add2[3]),.Cout(carry2[4]));
  multBlock mult25(.x(A[5]),.y(add1[5]),.alt(B[2]),.Cin(carry2[4]),.S(add2[4]),.Cout(carry2[5]));
  multBlock mult26(.x(A[6]),.y(add1[6]),.alt(B[2]),.Cin(carry2[5]),.S(add2[5]),.Cout(carry2[6]));
  multBlock mult27(.x(A[7]),.y(add1[7]),.alt(B[2]),.Cin(carry2[6]),.S(add2[6]),.Cout(carry2[7]));
  multBlock mult28(.x(A[8]),.y(add1[8]),.alt(B[2]),.Cin(carry2[7]),.S(add2[7]),.Cout(carry2[8]));
  multBlock mult29(.x(A[9]),.y(add1[9]),.alt(B[2]),.Cin(carry2[8]),.S(add2[8]),.Cout(carry2[9]));
  multBlock mult210(.x(A[10]),.y(add1[10]),.alt(B[2]),.Cin(carry2[9]),.S(add2[9]),.Cout(carry2[10]));
  multBlock mult211(.x(A[11]),.y(add1[11]),.alt(B[2]),.Cin(carry2[10]),.S(add2[10]),.Cout(carry2[11]));
  multBlock mult212(.x(A[12]),.y(add1[12]),.alt(B[2]),.Cin(carry2[11]),.S(add2[11]),.Cout(carry2[12]));
  multBlock mult213(.x(A[13]),.y(add1[13]),.alt(B[2]),.Cin(carry2[12]),.S(add2[12]),.Cout(carry2[13]));
  multBlock mult214(.x(A[14]),.y(add1[14]),.alt(B[2]),.Cin(carry2[13]),.S(add2[13]),.Cout(carry2[14]));
  multBlock mult215(.x(A[15]),.y(carry1[15]),.alt(B[2]),.Cin(carry2[14]),.S(add2[14]),.Cout(carry2[15]));
  //4th row of multiplier blocks
  multBlock mult30(.x(A[0]),.y(add2[0]),.alt(B[3]),.Cin(zero),.S(result[3]),.Cout(carry3[0]));
  multBlock mult31(.x(A[1]),.y(add2[1]),.alt(B[3]),.Cin(carry3[0]),.S(add3[0]),.Cout(carry3[1]));
  multBlock mult32(.x(A[2]),.y(add2[2]),.alt(B[3]),.Cin(carry3[1]),.S(add3[1]),.Cout(carry3[2]));
  multBlock mult33(.x(A[3]),.y(add2[3]),.alt(B[3]),.Cin(carry3[2]),.S(add3[2]),.Cout(carry3[3]));
  multBlock mult34(.x(A[4]),.y(add2[4]),.alt(B[3]),.Cin(carry3[3]),.S(add3[3]),.Cout(carry3[4]));
  multBlock mult35(.x(A[5]),.y(add2[5]),.alt(B[3]),.Cin(carry3[4]),.S(add3[4]),.Cout(carry3[5]));
  multBlock mult36(.x(A[6]),.y(add2[6]),.alt(B[3]),.Cin(carry3[5]),.S(add3[5]),.Cout(carry3[6]));
  multBlock mult37(.x(A[7]),.y(add2[7]),.alt(B[3]),.Cin(carry3[6]),.S(add3[6]),.Cout(carry3[7]));
  multBlock mult38(.x(A[8]),.y(add2[8]),.alt(B[3]),.Cin(carry3[7]),.S(add3[7]),.Cout(carry3[8]));
  multBlock mult39(.x(A[9]),.y(add2[9]),.alt(B[3]),.Cin(carry3[8]),.S(add3[8]),.Cout(carry3[9]));
  multBlock mult310(.x(A[10]),.y(add2[10]),.alt(B[3]),.Cin(carry3[9]),.S(add3[9]),.Cout(carry3[10]));
  multBlock mult311(.x(A[11]),.y(add2[11]),.alt(B[3]),.Cin(carry3[10]),.S(add3[10]),.Cout(carry3[11]));
  multBlock mult312(.x(A[12]),.y(add2[12]),.alt(B[3]),.Cin(carry3[11]),.S(add3[11]),.Cout(carry3[12]));
  multBlock mult313(.x(A[13]),.y(add2[13]),.alt(B[3]),.Cin(carry3[12]),.S(add3[12]),.Cout(carry3[13]));
  multBlock mult314(.x(A[14]),.y(add2[14]),.alt(B[3]),.Cin(carry3[13]),.S(add3[13]),.Cout(carry3[14]));
  multBlock mult315(.x(A[15]),.y(carry2[15]),.alt(B[3]),.Cin(carry3[14]),.S(add3[14]),.Cout(carry3[15]));
  //5th row of multiplier blocks
  multBlock mult40(.x(A[0]),.y(add3[0]),.alt(B[4]),.Cin(zero),.S(result[4]),.Cout(carry4[0]));
  multBlock mult41(.x(A[1]),.y(add3[1]),.alt(B[4]),.Cin(carry4[0]),.S(add4[0]),.Cout(carry4[1]));
  multBlock mult42(.x(A[2]),.y(add3[2]),.alt(B[4]),.Cin(carry4[1]),.S(add4[1]),.Cout(carry4[2]));
  multBlock mult43(.x(A[3]),.y(add3[3]),.alt(B[4]),.Cin(carry4[2]),.S(add4[2]),.Cout(carry4[3]));
  multBlock mult44(.x(A[4]),.y(add3[4]),.alt(B[4]),.Cin(carry4[3]),.S(add4[3]),.Cout(carry4[4]));
  multBlock mult45(.x(A[5]),.y(add3[5]),.alt(B[4]),.Cin(carry4[4]),.S(add4[4]),.Cout(carry4[5]));
  multBlock mult46(.x(A[6]),.y(add3[6]),.alt(B[4]),.Cin(carry4[5]),.S(add4[5]),.Cout(carry4[6]));
  multBlock mult47(.x(A[7]),.y(add3[7]),.alt(B[4]),.Cin(carry4[6]),.S(add4[6]),.Cout(carry4[7]));
  multBlock mult48(.x(A[8]),.y(add3[8]),.alt(B[4]),.Cin(carry4[7]),.S(add4[7]),.Cout(carry4[8]));
  multBlock mult49(.x(A[9]),.y(add3[9]),.alt(B[4]),.Cin(carry4[8]),.S(add4[8]),.Cout(carry4[9]));
  multBlock mult410(.x(A[10]),.y(add3[10]),.alt(B[4]),.Cin(carry4[9]),.S(add4[9]),.Cout(carry4[10]));
  multBlock mult411(.x(A[11]),.y(add3[11]),.alt(B[4]),.Cin(carry4[10]),.S(add4[10]),.Cout(carry4[11]));
  multBlock mult412(.x(A[12]),.y(add3[12]),.alt(B[4]),.Cin(carry4[11]),.S(add4[11]),.Cout(carry4[12]));
  multBlock mult413(.x(A[13]),.y(add3[13]),.alt(B[4]),.Cin(carry4[12]),.S(add4[12]),.Cout(carry4[13]));
  multBlock mult414(.x(A[14]),.y(add3[14]),.alt(B[4]),.Cin(carry4[13]),.S(add4[13]),.Cout(carry4[14]));
  multBlock mult415(.x(A[15]),.y(carry3[15]),.alt(B[4]),.Cin(carry4[14]),.S(add4[14]),.Cout(carry4[15]));
  //6th row of multiplier blocks
  multBlock mult50(.x(A[0]),.y(add4[0]),.alt(B[5]),.Cin(zero),.S(result[5]),.Cout(carry5[0]));
  multBlock mult51(.x(A[1]),.y(add4[1]),.alt(B[5]),.Cin(carry5[0]),.S(add5[0]),.Cout(carry5[1]));
  multBlock mult52(.x(A[2]),.y(add4[2]),.alt(B[5]),.Cin(carry5[1]),.S(add5[1]),.Cout(carry5[2]));
  multBlock mult53(.x(A[3]),.y(add4[3]),.alt(B[5]),.Cin(carry5[2]),.S(add5[2]),.Cout(carry5[3]));
  multBlock mult54(.x(A[4]),.y(add4[4]),.alt(B[5]),.Cin(carry5[3]),.S(add5[3]),.Cout(carry5[4]));
  multBlock mult55(.x(A[5]),.y(add4[5]),.alt(B[5]),.Cin(carry5[4]),.S(add5[4]),.Cout(carry5[5]));
  multBlock mult56(.x(A[6]),.y(add4[6]),.alt(B[5]),.Cin(carry5[5]),.S(add5[5]),.Cout(carry5[6]));
  multBlock mult57(.x(A[7]),.y(add4[7]),.alt(B[5]),.Cin(carry5[6]),.S(add5[6]),.Cout(carry5[7]));
  multBlock mult58(.x(A[8]),.y(add4[8]),.alt(B[5]),.Cin(carry5[7]),.S(add5[7]),.Cout(carry5[8]));
  multBlock mult59(.x(A[9]),.y(add4[9]),.alt(B[5]),.Cin(carry5[8]),.S(add5[8]),.Cout(carry5[9]));
  multBlock mult510(.x(A[10]),.y(add4[10]),.alt(B[5]),.Cin(carry5[9]),.S(add5[9]),.Cout(carry5[10]));
  multBlock mult511(.x(A[11]),.y(add4[11]),.alt(B[5]),.Cin(carry5[10]),.S(add5[10]),.Cout(carry5[11]));
  multBlock mult512(.x(A[12]),.y(add4[12]),.alt(B[5]),.Cin(carry5[11]),.S(add5[11]),.Cout(carry5[12]));
  multBlock mult513(.x(A[13]),.y(add4[13]),.alt(B[5]),.Cin(carry5[12]),.S(add5[12]),.Cout(carry5[13]));
  multBlock mult514(.x(A[14]),.y(add4[14]),.alt(B[5]),.Cin(carry5[13]),.S(add5[13]),.Cout(carry5[14]));
  multBlock mult515(.x(A[15]),.y(carry4[15]),.alt(B[5]),.Cin(carry5[14]),.S(add5[14]),.Cout(carry5[15]));
  //7th row of multiplier blocks
  multBlock mult60(.x(A[0]),.y(add5[0]),.alt(B[6]),.Cin(zero),.S(result[6]),.Cout(carry6[0]));
  multBlock mult61(.x(A[1]),.y(add5[1]),.alt(B[6]),.Cin(carry6[0]),.S(add6[0]),.Cout(carry6[1]));
  multBlock mult62(.x(A[2]),.y(add5[2]),.alt(B[6]),.Cin(carry6[1]),.S(add6[1]),.Cout(carry6[2]));
  multBlock mult63(.x(A[3]),.y(add5[3]),.alt(B[6]),.Cin(carry6[2]),.S(add6[2]),.Cout(carry6[3]));
  multBlock mult64(.x(A[4]),.y(add5[4]),.alt(B[6]),.Cin(carry6[3]),.S(add6[3]),.Cout(carry6[4]));
  multBlock mult65(.x(A[5]),.y(add5[5]),.alt(B[6]),.Cin(carry6[4]),.S(add6[4]),.Cout(carry6[5]));
  multBlock mult66(.x(A[6]),.y(add5[6]),.alt(B[6]),.Cin(carry6[5]),.S(add6[5]),.Cout(carry6[6]));
  multBlock mult67(.x(A[7]),.y(add5[7]),.alt(B[6]),.Cin(carry6[6]),.S(add6[6]),.Cout(carry6[7]));
  multBlock mult68(.x(A[8]),.y(add5[8]),.alt(B[6]),.Cin(carry6[7]),.S(add6[7]),.Cout(carry6[8]));
  multBlock mult69(.x(A[9]),.y(add5[9]),.alt(B[6]),.Cin(carry6[8]),.S(add6[8]),.Cout(carry6[9]));
  multBlock mult610(.x(A[10]),.y(add5[10]),.alt(B[6]),.Cin(carry6[9]),.S(add6[9]),.Cout(carry6[10]));
  multBlock mult611(.x(A[11]),.y(add5[11]),.alt(B[6]),.Cin(carry6[10]),.S(add6[10]),.Cout(carry6[11]));
  multBlock mult612(.x(A[12]),.y(add5[12]),.alt(B[6]),.Cin(carry6[11]),.S(add6[11]),.Cout(carry6[12]));
  multBlock mult613(.x(A[13]),.y(add5[13]),.alt(B[6]),.Cin(carry6[12]),.S(add6[12]),.Cout(carry6[13]));
  multBlock mult614(.x(A[14]),.y(add5[14]),.alt(B[6]),.Cin(carry6[13]),.S(add6[13]),.Cout(carry6[14]));
  multBlock mult615(.x(A[15]),.y(add5[15]),.alt(B[6]),.Cin(carry6[14]),.S(add6[14]),.Cout(carry6[15]));
  //8th row of multiplier blocks
  multBlock mult70(.x(A[0]),.y(add6[0]),.alt(B[7]),.Cin(zero),.S(result[7]),.Cout(carry7[0]));
  multBlock mult71(.x(A[1]),.y(add6[1]),.alt(B[7]),.Cin(carry7[0]),.S(add7[0]),.Cout(carry7[1]));
  multBlock mult72(.x(A[2]),.y(add6[2]),.alt(B[7]),.Cin(carry7[1]),.S(add7[1]),.Cout(carry7[2]));
  multBlock mult73(.x(A[3]),.y(add6[3]),.alt(B[7]),.Cin(carry7[2]),.S(add7[2]),.Cout(carry7[3]));
  multBlock mult74(.x(A[4]),.y(add6[4]),.alt(B[7]),.Cin(carry7[3]),.S(add7[3]),.Cout(carry7[4]));
  multBlock mult75(.x(A[5]),.y(add6[5]),.alt(B[7]),.Cin(carry7[4]),.S(add7[4]),.Cout(carry7[5]));
  multBlock mult76(.x(A[6]),.y(add6[6]),.alt(B[7]),.Cin(carry7[5]),.S(add7[5]),.Cout(carry7[6]));
  multBlock mult77(.x(A[7]),.y(add6[7]),.alt(B[7]),.Cin(carry7[6]),.S(add7[6]),.Cout(carry7[7]));
  multBlock mult78(.x(A[8]),.y(add6[8]),.alt(B[7]),.Cin(carry7[7]),.S(add7[7]),.Cout(carry7[8]));
  multBlock mult79(.x(A[9]),.y(add6[9]),.alt(B[7]),.Cin(carry7[8]),.S(add7[8]),.Cout(carry7[9]));
  multBlock mult710(.x(A[10]),.y(add6[10]),.alt(B[7]),.Cin(carry7[9]),.S(add7[9]),.Cout(carry7[10]));
  multBlock mult711(.x(A[11]),.y(add6[11]),.alt(B[7]),.Cin(carry7[10]),.S(add7[10]),.Cout(carry7[11]));
  multBlock mult712(.x(A[12]),.y(add6[12]),.alt(B[7]),.Cin(carry7[11]),.S(add7[11]),.Cout(carry7[12]));
  multBlock mult713(.x(A[13]),.y(add6[13]),.alt(B[7]),.Cin(carry7[12]),.S(add7[12]),.Cout(carry7[13]));
  multBlock mult714(.x(A[14]),.y(add6[14]),.alt(B[7]),.Cin(carry7[13]),.S(add7[13]),.Cout(carry7[14]));
  multBlock mult715(.x(A[15]),.y(add6[15]),.alt(B[7]),.Cin(carry7[14]),.S(add7[14]),.Cout(carry7[15]));
  //9th row of multiplier blocks
  multBlock mult80(.x(A[0]),.y(add7[0]),.alt(B[8]),.Cin(zero),.S(result[8]),.Cout(carry8[0]));
  multBlock mult81(.x(A[1]),.y(add7[1]),.alt(B[8]),.Cin(carry8[0]),.S(add8[0]),.Cout(carry8[1]));
  multBlock mult82(.x(A[2]),.y(add7[2]),.alt(B[8]),.Cin(carry8[1]),.S(add8[1]),.Cout(carry8[2]));
  multBlock mult83(.x(A[3]),.y(add7[3]),.alt(B[8]),.Cin(carry8[2]),.S(add8[2]),.Cout(carry8[3]));
  multBlock mult84(.x(A[4]),.y(add7[4]),.alt(B[8]),.Cin(carry8[3]),.S(add8[3]),.Cout(carry8[4]));
  multBlock mult85(.x(A[5]),.y(add7[5]),.alt(B[8]),.Cin(carry8[4]),.S(add8[4]),.Cout(carry8[5]));
  multBlock mult86(.x(A[6]),.y(add7[6]),.alt(B[8]),.Cin(carry8[5]),.S(add8[5]),.Cout(carry8[6]));
  multBlock mult87(.x(A[7]),.y(add7[7]),.alt(B[8]),.Cin(carry8[6]),.S(add8[6]),.Cout(carry8[7]));
  multBlock mult88(.x(A[8]),.y(add7[8]),.alt(B[8]),.Cin(carry8[7]),.S(add8[7]),.Cout(carry8[8]));
  multBlock mult89(.x(A[9]),.y(add7[9]),.alt(B[8]),.Cin(carry8[8]),.S(add8[8]),.Cout(carry8[9]));
  multBlock mult810(.x(A[10]),.y(add7[10]),.alt(B[8]),.Cin(carry8[9]),.S(add8[9]),.Cout(carry8[10]));
  multBlock mult811(.x(A[11]),.y(add7[11]),.alt(B[8]),.Cin(carry8[10]),.S(add8[10]),.Cout(carry8[11]));
  multBlock mult812(.x(A[12]),.y(add7[12]),.alt(B[8]),.Cin(carry8[11]),.S(add8[11]),.Cout(carry8[12]));
  multBlock mult813(.x(A[13]),.y(add7[13]),.alt(B[8]),.Cin(carry8[12]),.S(add8[12]),.Cout(carry8[13]));
  multBlock mult814(.x(A[14]),.y(add7[14]),.alt(B[8]),.Cin(carry8[13]),.S(add8[13]),.Cout(carry8[14]));
  multBlock mult815(.x(A[15]),.y(add7[15]),.alt(B[8]),.Cin(carry8[14]),.S(add8[14]),.Cout(carry8[15]));
  //10th row of multiplier blocks
  multBlock mult90(.x(A[0]),.y(add8[0]),.alt(B[9]),.Cin(zero),.S(result[9]),.Cout(carry9[0]));
  multBlock mult91(.x(A[1]),.y(add8[1]),.alt(B[9]),.Cin(carry9[0]),.S(add9[0]),.Cout(carry9[1]));
  multBlock mult92(.x(A[2]),.y(add8[2]),.alt(B[9]),.Cin(carry9[1]),.S(add9[1]),.Cout(carry9[2]));
  multBlock mult93(.x(A[3]),.y(add8[3]),.alt(B[9]),.Cin(carry9[2]),.S(add9[2]),.Cout(carry9[3]));
  multBlock mult94(.x(A[4]),.y(add8[4]),.alt(B[9]),.Cin(carry9[3]),.S(add9[3]),.Cout(carry9[4]));
  multBlock mult95(.x(A[5]),.y(add8[5]),.alt(B[9]),.Cin(carry9[4]),.S(add9[4]),.Cout(carry9[5]));
  multBlock mult96(.x(A[6]),.y(add8[6]),.alt(B[9]),.Cin(carry9[5]),.S(add9[5]),.Cout(carry9[6]));
  multBlock mult97(.x(A[7]),.y(add8[7]),.alt(B[9]),.Cin(carry9[6]),.S(add9[6]),.Cout(carry9[7]));
  multBlock mult98(.x(A[8]),.y(add8[8]),.alt(B[9]),.Cin(carry9[7]),.S(add9[7]),.Cout(carry9[8]));
  multBlock mult99(.x(A[9]),.y(add8[9]),.alt(B[9]),.Cin(carry9[8]),.S(add9[8]),.Cout(carry9[9]));
  multBlock mult910(.x(A[10]),.y(add8[10]),.alt(B[9]),.Cin(carry9[9]),.S(add9[9]),.Cout(carry9[10]));
  multBlock mult911(.x(A[11]),.y(add8[11]),.alt(B[9]),.Cin(carry9[10]),.S(add9[10]),.Cout(carry9[11]));
  multBlock mult912(.x(A[12]),.y(add8[12]),.alt(B[9]),.Cin(carry9[11]),.S(add9[11]),.Cout(carry9[12]));
  multBlock mult913(.x(A[13]),.y(add8[13]),.alt(B[9]),.Cin(carry9[12]),.S(add9[12]),.Cout(carry9[13]));
  multBlock mult914(.x(A[14]),.y(add8[14]),.alt(B[9]),.Cin(carry9[13]),.S(add9[13]),.Cout(carry9[14]));
  multBlock mult915(.x(A[15]),.y(add8[15]),.alt(B[9]),.Cin(carry9[14]),.S(add9[14]),.Cout(carry9[15]));
  //11th row of multiplier blocks
  multBlock mult100(.x(A[0]),.y(add9[0]),.alt(B[10]),.Cin(zero),.S(result[10]),.Cout(carry10[0]));
  multBlock mult101(.x(A[1]),.y(add9[1]),.alt(B[10]),.Cin(carry10[0]),.S(add10[0]),.Cout(carry10[1]));
  multBlock mult102(.x(A[2]),.y(add9[2]),.alt(B[10]),.Cin(carry10[1]),.S(add10[1]),.Cout(carry10[2]));
  multBlock mult103(.x(A[3]),.y(add9[3]),.alt(B[10]),.Cin(carry10[2]),.S(add10[2]),.Cout(carry10[3]));
  multBlock mult104(.x(A[4]),.y(add9[4]),.alt(B[10]),.Cin(carry10[3]),.S(add10[3]),.Cout(carry10[4]));
  multBlock mult105(.x(A[5]),.y(add9[5]),.alt(B[10]),.Cin(carry10[4]),.S(add10[4]),.Cout(carry10[5]));
  multBlock mult106(.x(A[6]),.y(add9[6]),.alt(B[10]),.Cin(carry10[5]),.S(add10[5]),.Cout(carry10[6]));
  multBlock mult107(.x(A[7]),.y(add9[7]),.alt(B[10]),.Cin(carry10[6]),.S(add10[6]),.Cout(carry10[7]));
  multBlock mult108(.x(A[8]),.y(add9[8]),.alt(B[10]),.Cin(carry10[7]),.S(add10[7]),.Cout(carry10[8]));
  multBlock mult109(.x(A[9]),.y(add9[9]),.alt(B[10]),.Cin(carry10[8]),.S(add10[8]),.Cout(carry10[9]));
  multBlock mult1010(.x(A[10]),.y(add9[10]),.alt(B[10]),.Cin(carry10[9]),.S(add10[9]),.Cout(carry10[10]));
  multBlock mult1011(.x(A[11]),.y(add9[11]),.alt(B[10]),.Cin(carry10[10]),.S(add10[10]),.Cout(carry10[11]));
  multBlock mult1012(.x(A[12]),.y(add9[12]),.alt(B[10]),.Cin(carry10[11]),.S(add10[11]),.Cout(carry10[12]));
  multBlock mult1013(.x(A[13]),.y(add9[13]),.alt(B[10]),.Cin(carry10[12]),.S(add10[12]),.Cout(carry10[13]));
  multBlock mult1014(.x(A[14]),.y(add9[14]),.alt(B[10]),.Cin(carry10[13]),.S(add10[13]),.Cout(carry10[14]));
  multBlock mult1015(.x(A[15]),.y(add9[15]),.alt(B[10]),.Cin(carry10[14]),.S(add10[14]),.Cout(carry10[15]));
  //12th row of multiplier blocks
  multBlock mult11_0(.x(A[0]),.y(add10[0]),.alt(B[11]),.Cin(zero),.S(result[11]),.Cout(carry11[0]));
  multBlock mult11_1(.x(A[1]),.y(add10[1]),.alt(B[11]),.Cin(carry11[0]),.S(add11[0]),.Cout(carry11[1]));
  multBlock mult11_2(.x(A[2]),.y(add10[2]),.alt(B[11]),.Cin(carry11[1]),.S(add11[1]),.Cout(carry11[2]));
  multBlock mult11_3(.x(A[3]),.y(add10[3]),.alt(B[11]),.Cin(carry11[2]),.S(add11[2]),.Cout(carry11[3]));
  multBlock mult11_4(.x(A[4]),.y(add10[4]),.alt(B[11]),.Cin(carry11[3]),.S(add11[3]),.Cout(carry11[4]));
  multBlock mult11_5(.x(A[5]),.y(add10[5]),.alt(B[11]),.Cin(carry11[4]),.S(add11[4]),.Cout(carry11[5]));
  multBlock mult11_6(.x(A[6]),.y(add10[6]),.alt(B[11]),.Cin(carry11[5]),.S(add11[5]),.Cout(carry11[6]));
  multBlock mult117(.x(A[7]),.y(add10[7]),.alt(B[11]),.Cin(carry11[6]),.S(add11[6]),.Cout(carry11[7]));
  multBlock mult118(.x(A[8]),.y(add10[8]),.alt(B[11]),.Cin(carry11[7]),.S(add11[7]),.Cout(carry11[8]));
  multBlock mult119(.x(A[9]),.y(add10[9]),.alt(B[11]),.Cin(carry11[8]),.S(add11[8]),.Cout(carry11[9]));
  multBlock mult1110(.x(A[10]),.y(add10[10]),.alt(B[11]),.Cin(carry11[9]),.S(add11[9]),.Cout(carry11[10]));
  multBlock mult1111(.x(A[11]),.y(add10[11]),.alt(B[11]),.Cin(carry11[10]),.S(add11[10]),.Cout(carry11[11]));
  multBlock mult1112(.x(A[12]),.y(add10[12]),.alt(B[11]),.Cin(carry11[11]),.S(add11[11]),.Cout(carry11[12]));
  multBlock mult1113(.x(A[13]),.y(add10[13]),.alt(B[11]),.Cin(carry11[12]),.S(add11[12]),.Cout(carry11[13]));
  multBlock mult1114(.x(A[14]),.y(add10[14]),.alt(B[11]),.Cin(carry11[13]),.S(add11[13]),.Cout(carry11[14]));
  multBlock mult1115(.x(A[15]),.y(add10[15]),.alt(B[11]),.Cin(carry11[14]),.S(add11[14]),.Cout(carry11[15]));
  //13th row of multiplier blocks
  multBlock mult120(.x(A[0]),.y(add11[0]),.alt(B[12]),.Cin(zero),.S(result[12]),.Cout(carry12[0]));
  multBlock mult121(.x(A[1]),.y(add11[1]),.alt(B[12]),.Cin(carry12[0]),.S(add12[0]),.Cout(carry12[1]));
  multBlock mult122(.x(A[2]),.y(add11[2]),.alt(B[12]),.Cin(carry12[1]),.S(add12[1]),.Cout(carry12[2]));
  multBlock mult123(.x(A[3]),.y(add11[3]),.alt(B[12]),.Cin(carry12[2]),.S(add12[2]),.Cout(carry12[3]));
  multBlock mult124(.x(A[4]),.y(add11[4]),.alt(B[12]),.Cin(carry12[3]),.S(add12[3]),.Cout(carry12[4]));
  multBlock mult125(.x(A[5]),.y(add11[5]),.alt(B[12]),.Cin(carry12[4]),.S(add12[4]),.Cout(carry12[5]));
  multBlock mult126(.x(A[6]),.y(add11[6]),.alt(B[12]),.Cin(carry12[5]),.S(add12[5]),.Cout(carry12[6]));
  multBlock mult127(.x(A[7]),.y(add11[7]),.alt(B[12]),.Cin(carry12[6]),.S(add12[6]),.Cout(carry12[7]));
  multBlock mult128(.x(A[8]),.y(add11[8]),.alt(B[12]),.Cin(carry12[7]),.S(add12[7]),.Cout(carry12[8]));
  multBlock mult129(.x(A[9]),.y(add11[9]),.alt(B[12]),.Cin(carry12[8]),.S(add12[8]),.Cout(carry12[9]));
  multBlock mult1210(.x(A[10]),.y(add11[10]),.alt(B[12]),.Cin(carry12[9]),.S(add12[9]),.Cout(carry12[10]));
  multBlock mult1211(.x(A[11]),.y(add11[11]),.alt(B[12]),.Cin(carry12[10]),.S(add12[10]),.Cout(carry12[11]));
  multBlock mult1212(.x(A[12]),.y(add11[12]),.alt(B[12]),.Cin(carry12[11]),.S(add12[11]),.Cout(carry12[12]));
  multBlock mult1213(.x(A[13]),.y(add11[13]),.alt(B[12]),.Cin(carry12[12]),.S(add12[12]),.Cout(carry12[13]));
  multBlock mult1214(.x(A[14]),.y(add11[14]),.alt(B[12]),.Cin(carry12[13]),.S(add12[13]),.Cout(carry12[14]));
  multBlock mult1215(.x(A[15]),.y(add11[15]),.alt(B[12]),.Cin(carry12[14]),.S(add12[14]),.Cout(carry12[15]));
  //14th row of multiplier blocks
  multBlock mult130(.x(A[0]),.y(add12[0]),.alt(B[13]),.Cin(zero),.S(result[13]),.Cout(carry13[0]));
  multBlock mult131(.x(A[1]),.y(add12[1]),.alt(B[13]),.Cin(carry13[0]),.S(add13[0]),.Cout(carry13[1]));
  multBlock mult132(.x(A[2]),.y(add12[2]),.alt(B[13]),.Cin(carry13[1]),.S(add13[1]),.Cout(carry13[2]));
  multBlock mult133(.x(A[3]),.y(add12[3]),.alt(B[13]),.Cin(carry13[2]),.S(add13[2]),.Cout(carry13[3]));
  multBlock mult134(.x(A[4]),.y(add12[4]),.alt(B[13]),.Cin(carry13[3]),.S(add13[3]),.Cout(carry13[4]));
  multBlock mult135(.x(A[5]),.y(add12[5]),.alt(B[13]),.Cin(carry13[4]),.S(add13[4]),.Cout(carry13[5]));
  multBlock mult136(.x(A[6]),.y(add12[6]),.alt(B[13]),.Cin(carry13[5]),.S(add13[5]),.Cout(carry13[6]));
  multBlock mult137(.x(A[7]),.y(add12[7]),.alt(B[13]),.Cin(carry13[6]),.S(add13[6]),.Cout(carry13[7]));
  multBlock mult138(.x(A[8]),.y(add12[8]),.alt(B[13]),.Cin(carry13[7]),.S(add13[7]),.Cout(carry13[8]));
  multBlock mult139(.x(A[9]),.y(add12[9]),.alt(B[13]),.Cin(carry13[8]),.S(add13[8]),.Cout(carry13[9]));
  multBlock mult1310(.x(A[10]),.y(add12[10]),.alt(B[13]),.Cin(carry13[9]),.S(add13[9]),.Cout(carry13[10]));
  multBlock mult1311(.x(A[11]),.y(add12[11]),.alt(B[13]),.Cin(carry13[10]),.S(add13[10]),.Cout(carry13[11]));
  multBlock mult1312(.x(A[12]),.y(add12[12]),.alt(B[13]),.Cin(carry13[11]),.S(add13[11]),.Cout(carry13[12]));
  multBlock mult1313(.x(A[13]),.y(add12[13]),.alt(B[13]),.Cin(carry13[12]),.S(add13[12]),.Cout(carry13[13]));
  multBlock mult1314(.x(A[14]),.y(add12[14]),.alt(B[13]),.Cin(carry13[13]),.S(add13[13]),.Cout(carry13[14]));
  multBlock mult1315(.x(A[15]),.y(add12[15]),.alt(B[13]),.Cin(carry13[14]),.S(add13[14]),.Cout(carry13[15]));
  //15th row of multiplier blocks
  multBlock mult140(.x(A[0]),.y(add13[0]),.alt(B[14]),.Cin(zero),.S(result[14]),.Cout(carry14[0]));
  multBlock mult141(.x(A[1]),.y(add13[1]),.alt(B[14]),.Cin(carry14[0]),.S(add14[0]),.Cout(carry14[1]));
  multBlock mult142(.x(A[2]),.y(add13[2]),.alt(B[14]),.Cin(carry14[1]),.S(add14[1]),.Cout(carry14[2]));
  multBlock mult143(.x(A[3]),.y(add13[3]),.alt(B[14]),.Cin(carry14[2]),.S(add14[2]),.Cout(carry14[3]));
  multBlock mult144(.x(A[4]),.y(add13[4]),.alt(B[14]),.Cin(carry14[3]),.S(add14[3]),.Cout(carry14[4]));
  multBlock mult145(.x(A[5]),.y(add13[5]),.alt(B[14]),.Cin(carry14[4]),.S(add14[4]),.Cout(carry14[5]));
  multBlock mult146(.x(A[6]),.y(add13[6]),.alt(B[14]),.Cin(carry14[5]),.S(add14[5]),.Cout(carry14[6]));
  multBlock mult147(.x(A[7]),.y(add13[7]),.alt(B[14]),.Cin(carry14[6]),.S(add14[6]),.Cout(carry14[7]));
  multBlock mult148(.x(A[8]),.y(add13[8]),.alt(B[14]),.Cin(carry14[7]),.S(add14[7]),.Cout(carry14[8]));
  multBlock mult149(.x(A[9]),.y(add13[9]),.alt(B[14]),.Cin(carry14[8]),.S(add14[8]),.Cout(carry14[9]));
  multBlock mult1410(.x(A[10]),.y(add13[10]),.alt(B[14]),.Cin(carry14[9]),.S(add14[9]),.Cout(carry14[10]));
  multBlock mult1411(.x(A[11]),.y(add13[11]),.alt(B[14]),.Cin(carry14[10]),.S(add14[10]),.Cout(carry14[11]));
  multBlock mult1412(.x(A[12]),.y(add13[12]),.alt(B[14]),.Cin(carry14[11]),.S(add14[11]),.Cout(carry14[12]));
  multBlock mult1413(.x(A[13]),.y(add13[13]),.alt(B[14]),.Cin(carry14[12]),.S(add14[12]),.Cout(carry14[13]));
  multBlock mult1414(.x(A[14]),.y(add13[14]),.alt(B[14]),.Cin(carry14[13]),.S(add14[13]),.Cout(carry14[14]));
  multBlock mult1415(.x(A[15]),.y(add13[15]),.alt(B[14]),.Cin(carry14[14]),.S(add14[14]),.Cout(carry14[15]));
  //16th row of multiplier blocks
  multBlock mult150(.x(A[0]),.y(add14[0]),.alt(B[15]),.Cin(zero),.S(result[15]),.Cout(carry15[0]));
  multBlock mult151(.x(A[1]),.y(add14[1]),.alt(B[15]),.Cin(carry15[0]),.S(result[16]),.Cout(carry15[1]));
  multBlock mult152(.x(A[2]),.y(add14[2]),.alt(B[15]),.Cin(carry15[1]),.S(result[17]),.Cout(carry15[2]));
  multBlock mult153(.x(A[3]),.y(add14[3]),.alt(B[15]),.Cin(carry15[2]),.S(result[18]),.Cout(carry15[3]));
  multBlock mult154(.x(A[4]),.y(add14[4]),.alt(B[15]),.Cin(carry15[3]),.S(result[19]),.Cout(carry15[4]));
  multBlock mult155(.x(A[5]),.y(add14[5]),.alt(B[15]),.Cin(carry15[4]),.S(result[20]),.Cout(carry15[5]));
  multBlock mult156(.x(A[6]),.y(add14[6]),.alt(B[15]),.Cin(carry15[5]),.S(result[21]),.Cout(carry15[6]));
  multBlock mult157(.x(A[7]),.y(add14[7]),.alt(B[15]),.Cin(carry15[6]),.S(result[22]),.Cout(carry15[7]));
  multBlock mult158(.x(A[8]),.y(add14[8]),.alt(B[15]),.Cin(carry15[7]),.S(result[23]),.Cout(carry15[8]));
  multBlock mult159(.x(A[9]),.y(add14[9]),.alt(B[15]),.Cin(carry15[8]),.S(result[24]),.Cout(carry15[9]));
  multBlock mult1510(.x(A[10]),.y(add14[10]),.alt(B[15]),.Cin(carry15[9]),.S(result[25]),.Cout(carry15[10]));
  multBlock mult1511(.x(A[11]),.y(add14[11]),.alt(B[15]),.Cin(carry15[10]),.S(result[26]),.Cout(carry15[11]));
  multBlock mult1512(.x(A[12]),.y(add14[12]),.alt(B[15]),.Cin(carry15[11]),.S(result[27]),.Cout(carry15[12]));
  multBlock mult1513(.x(A[13]),.y(add14[13]),.alt(B[15]),.Cin(carry15[12]),.S(result[28]),.Cout(carry15[13]));
  multBlock mult1514(.x(A[14]),.y(add14[14]),.alt(B[15]),.Cin(carry15[13]),.S(result[29]),.Cout(carry15[14]));
  multBlock mult1515(.x(A[15]),.y(add14[15]),.alt(B[15]),.Cin(carry15[14]),.S(result[30]),.Cout(result[31]));
  initial begin
    $display("%b",result);
    $finish;
  end
endmodule
